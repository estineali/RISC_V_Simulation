module RegisterFile
(
	input [4:0] rs1, rs2, rd,
	input [63:0] WriteData,
	input clk, reset, RegWrite,
	output reg [63:0] ReadData1, ReadData2
);

	reg [63:0] Registers [31:0];
	initial
	begin
		Registers[0] <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
		Registers[1] <= 64'b1001011000101111011000100001110110011001100101110101000000011011;
		Registers[2] <= 64'b1000111011111110000010111011001110100100100001010010100000010010;
		Registers[3] <= 64'b1001110110000101111010110010001110101011110101110000111000011110;
		Registers[4] <= 64'b1001001111000011011000001001110110110010011001111110110111000010;
		Registers[5] <= 64'b1011011110011100110101100100111010110101110101010101111001111110;
		Registers[6] <= 64'b1111011110100011100011010101000000010000100000110111101110100000;
		Registers[7] <= 64'b1001000000000010100000001100110110001001101110100010100111011011;
		Registers[8] <= 64'b0011010101100101100110000010111000101111011101111110110010000101;
		Registers[9] <= 64'b1000101010101101001000101101001001101111010111000010101010111010;
		Registers[10] <= 64'b1101001101010001011010010000100101110001001100000110011100000001;
		Registers[11] <= 64'b0010100110110101000011100001000110100011111001111000101001101010;
		Registers[12] <= 64'b1111111010101110000001110111010101100011000110100110111111100111;
		Registers[13] <= 64'b1110110000111110010100000100111000101100111010100111011111101000;
		Registers[14] <= 64'b1100110001110000001000010110010011101001111011001011011110111011;
		Registers[15] <= 64'b0101000111010111001011001010001011111001110001100000111011000101;
		Registers[16] <= 64'b0001100110100100101101001001101011001110010100100010111001110010;
		Registers[17] <= 64'b1000101011000001111011100000011010010111101101000010010101100000;
		Registers[18] <= 64'b0101011100110000110101000011000000001011111011100101010011010111;
		Registers[19] <= 64'b0111100011001100000010001001100100001110101011110001100001111110;
		Registers[20] <= 64'b0011010100100100101110001101111101000010010000101000001101110101;
		Registers[21] <= 64'b0000111110011110000000011100101111010110100011011010010111011111;
		Registers[22] <= 64'b0111011100110000000010001011011111100101010100111001111110000111;
		Registers[23] <= 64'b0010011101110100010010011001010001101010101000101101111001011101;
		Registers[24] <= 64'b0100110000111000010100101110001001010110111100011011111110100101;
		Registers[25] <= 64'b0101000101000100001101111110011100001010010100011010100001010110;
		Registers[26] <= 64'b0110000001101100000000100001001011101110001101011100001100011000;
		Registers[27] <= 64'b1101010101100111001110001101101101001111000110011010110100000000;
		Registers[28] <= 64'b0011111000101000100001010111110100000011000010011110001011011010;
		Registers[29] <= 64'b0111000000001011001001011101001001010110011010010001110101110100;
		Registers[30] <= 64'b1101010111001001111000000011100011011101111010011010101011110110;
		Registers[31] <= 64'b1001111101011010001010101001101100101111111011100100100010011110;
	end

	//Writing Data
	always @ (posedge clk)
	begin
		if (RegWrite == 1'b1)
			Registers[rd] = WriteData;
	end

	//Reseting ReadData ports
	always @ (reset)
	begin
		ReadData1 = 64'b0;
		ReadData2 = 64'b0; 
	end

	//output Data in ReadData Ports 
	always @ (rs1 or rs2 or reset)
	begin
		ReadData1 = Registers [rs1];
		ReadData2 = Registers [rs2];
	end

endmodule